module main

import echo


fn main(){
	mut e := echo.new_echo()

	e.run(8888)
}