module echo
//
// pub fn init_state() fn {
//
// 	mut state := 0
//
// 	return fn(){
//
// 	}
// }

// generic is not yet